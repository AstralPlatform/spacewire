// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51

module spacewire (
  input logic clk_i,
  input logic rst_ni
);

endmodule: spacewire
