library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;

library work;
use work.records_pkg.all;
use work.segm_mips_const_pkg.all;

entity spacewire is port(
  clk_i	 : in STD_LOGIC;
  rst_ni : in STD_LOGIC;
);
end spacewire;

architecture spacewire_arc of spacewire is

end spacewire_arc;
